* Current measure

.MODEL D1N4148 D (IS=4.352E-9 N=1.906 BV=110 IBV=0.0001 RS=0.6458 CJO=7.048E-13 VJ=0.869 M=0.03 FC=0.5 TT=3.48E-9 )


I1 1 0 AC 0 DC 0 PULSE( 0 65mA 0 1uS 1uS 150uS 1.6mS ) 
I2 1 0 AC 0 DC 0 PULSE( 0 -65mA 152uS 1uS 1uS 150uS 1.6mS ) 
R1 1 0 90.9R 
D1 1 2 D1N4148
D2 0 2 D1N4148
D3 3 1 D1N4148
D4 3 0 D1N4148
R2 2 3 475K
C1 2 3 1000uF

